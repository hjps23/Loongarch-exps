`timescale 1ns / 1ps
module redirect_unit(
    // ID�׶���Ϣ
    input  wire [4:0]  rj_in,
    input  wire [4:0]  rkd_in,
    // EX�׶���Ϣ
    input  wire        ex_gr_we,
    input  wire [4:0]  ex_dest,
    
    // MEM�׶���Ϣ  
    input  wire        mem_gr_we,
    input  wire [4:0]  mem_dest,
    
    // WB�׶���Ϣ
    input  wire        wb_gr_we,
    input  wire [4:0]  wb_dest,
    
    // �ض�������ź�
    output reg  [1:0]  rj_redirect,
    output reg  [1:0]  rkd_redirect
);


// rj�ض����߼�
always @(*) begin
    if (ex_gr_we && ex_dest != 5'b0 && ex_dest == rj_in) begin
        rj_redirect = 2'b01;  // ��EX�׶��ض���
    end else if ((mem_gr_we && mem_dest != 5'b0 && mem_dest == rj_in)) begin
        rj_redirect = 2'b10;  // ��MEM�׶��ض���
    end else if (wb_gr_we && wb_dest != 5'b0 && wb_dest == rj_in) begin
        rj_redirect = 2'b11;  // ��WB�׶��ض���
    end else begin
        rj_redirect = 2'b00;  // ���ض���
    end
end

// rk/rd�ض����߼�
always @(*) begin
    if (ex_gr_we && ex_dest != 5'b0 && ex_dest == rkd_in) begin
        rkd_redirect = 2'b01;  // ��EX�׶��ض���
    end else if ((mem_gr_we && mem_dest != 5'b0 && mem_dest == rkd_in)) begin
        rkd_redirect = 2'b10;  // ��MEM�׶��ض���
    end else if (wb_gr_we && wb_dest != 5'b0 && wb_dest == rkd_in) begin
        rkd_redirect = 2'b11;  // ��WB�׶��ض���
    end else begin
        rkd_redirect = 2'b00;  // ���ض���
    end
end

endmodule